use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(31 downto 0));
end uMem;

architecture Behavioral of uMem is

-- TODO: understand what is going on here

-- micro Memory
type u_mem_t is array (0 to 17) of unsigned(31 downto 0);
constant u_mem_c : u_mem_t :=
   -- NaN  ALU   TB   FB S P LC  SEQ    uAddr
  (b"0000_0000_0111_0011_0_0_00_0000_00000000", -- ASR:=PC
   b"0000_0000_0010_0001_0_1_00_0000_00000000", -- IR:=PM, PC:=PC+1
   b"0000_0000_0000_0000_0_0_00_0010_00000000", -- uPC := K2
   b"0000_0000_0000_0000_0_0_00_0000_00000000", -- 
   b"0000_0100_0111_0000_0_0_00_0000_00000000", -- 
   b"0000_0100_0111_0000_0_0_00_0000_00000000", -- 
   b"0000_0100_0111_0000_0_1_00_0000_00000000", -- 
   b"0000_1000_0111_0000_0_0_00_0000_00000000", -- 
   b"0000_0101_0111_0000_0_0_00_0000_00000000", -- 
   b"0000_1011_0000_0000_0_0_00_0000_00000000", -- 
   b"0000_1011_0000_0000_0_0_00_0000_00000000",
   b"0000_1010_0000_0000_0_0_00_0000_00000000",
   b"0000_0000_0000_0000_0_0_00_0000_00000000",
   b"0000_0000_0000_0000_0_0_00_0000_00000000",
   b"0000_0000_0000_0000_0_0_00_0000_00000000",
   b"0000_0000_0000_0000_0_0_00_0000_00000000",
   b"0000_0000_0000_0000_0_0_00_0000_00000000",
   b"0000_0000_0000_0000_0_0_00_0000_00000000");

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
