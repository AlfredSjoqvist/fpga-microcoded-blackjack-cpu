library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(7 downto 0);
    uData : out unsigned(31 downto 0));
end uMem;

architecture Behavioral of uMem is

-- TODO: understand what is going on here

-- micro Memory
type u_mem_t is array (0 to 255) of unsigned(31 downto 0);
constant u_mem_c : u_mem_t :=
   -- NaN  ALU   TB   FB GrPcLc  SEQ    uAddr
  (b"0000_0000_0111_0011_0_0_00_0000_00000000", -- ASR:=PC
   b"0000_0000_0010_0001_0_1_00_0000_00000000", -- IR  := PM, PC:=PC+1
   b"0000_0000_0000_0000_0_0_00_0010_00000000", -- uPC := K2
   b"0000_0000_0000_0000_0_0_00_0001_00000000", -- uPC := K1               ; Immediate/Implicit
   b"0000_0000_0001_0011_0_0_00_0001_00000000", -- ASR := IR, uPC := K1    ;   Direct
   b"0000_0000_0001_0011_0_0_00_0000_00000000", -- ASR := IR               ; Indirect                 
   b"0000_0000_0010_0011_0_0_00_0001_00000000", -- ASR := PM, uPC := K1    ; 
   b"0000_0001_0001_0000_0_0_00_0000_00000000", -- AR  := IR               ; Indexed
   b"0001_0100_0110_0000_1_0_00_0000_00000000", -- AR  := GrX+AR (noflag), GrSu = 1 ;
   b"0000_0000_0100_0011_0_0_00_0001_00000000", -- ASR := AR, uPC = K1     ;
   b"0000_0001_0111_0000_0_0_00_0000_00000000", -- AR := PC                ; Relative
   b"0001_0100_0001_0000_0_0_00_0000_00000000", -- AR := IR+AR (noflag)    ;
   b"0000_0000_0100_0111_0_0_00_0001_00000000", -- ASR := AR, uPC = K1     ;
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   
   b"0000_0000_0010_0110_0_0_00_0011_00000000", -- #LD   (mode, grx, adr)  ; GrX := PM(adr), uPC := 0
   b"0000_0000_0110_0010_0_0_00_0011_00000000", -- #ST   (mode, grx, adr)  ; PM(adr) := GrX, uPC := 0
   b"0000_0001_0000_0000_0_0_00_0000_00000000", -- #CMP  (mode, grx, adr)  ; AR := GrX
   b"0000_0101_0010_0000_0_0_00_0011_00000000", --                         ; AR := PM(adr) - AR, uPC := 0
   b"0000_0001_0110_0000_0_0_00_0000_00000000", -- #ADD  (mode, grx, adr)  ; AR  := GrX
   b"0000_0100_0010_0000_0_0_00_0000_00000000", --                         ; AR  := PM(adr) + AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0 
   b"0000_0001_0110_0000_0_0_00_0000_00000000", -- #SUB  (mode, grx, adr)  ; AR := GrX
   b"0000_0101_0010_0000_0_0_00_0000_00000000", --                         ; AR := PM(adr) - AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0
   b"0000_0001_0110_0000_0_0_00_0000_00000000", -- #AND  (mode, grx, adr)  ; AR := GrX
   b"0000_0110_0010_0000_0_0_00_0000_00000000", --                         ; AR := PM(adr) AND AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0
   b"0000_0001_0110_0000_0_0_00_0000_00000000", -- #OR   (mode, grx, adr)  ; AR := GrX
   b"0000_0111_0010_0000_0_0_00_0000_00000000", --                         ; AR := PM(adr) OR AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0

   b"0000_0001_0110_0000_0_0_00_0000_00000000", -- #MUL  (mode, grx, adr)  ; AR := GrX
   b"0000_1000_0010_0000_0_0_00_0000_00000000", --                         ; AR := PM(adr) * AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0
   b"0000_0001_0110_0000_0_0_00_0000_00000000", -- #MULS (mode, grx, adr)  ; AR := GrX
   b"0000_1001_0010_0000_0_0_00_0000_00000000", --                         ; AR := PM(adr) *(signed) AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0
   b"0000_0001_0010_0000_0_0_00_0000_00000000", -- #LSR  (mode, grx, adr)  ; AR := PM(adr)
   b"0000_1010_0000_0000_0_0_00_0000_00000000", --                         ; AR := lsr AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0
   b"0000_0001_0010_0000_0_0_00_0000_00000000", -- #LSL  (mode, grx, adr)  ; AR := PM(adr)
   b"0000_1011_0000_0000_0_0_00_0000_00000000", --                         ; AR := lsl AR
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0
   b"0000_0010_0010_0000_0_0_00_0000_00000000", -- #INV  (mode, grx, adr)  ; AR  := -PM(adr)
   b"0000_0000_0100_0110_0_0_00_0011_00000000", --                         ; GrX := AR, uPC := 0 
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --                         
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_1111_00000000", -- #HALT (----, ---, ---)  ; HALT

   b"0000_0000_0000_0000_0_0_00_0011_00000000", -- #JMP  (mode, ---, adr)  ; PC := PM(adr), uPC := 0
   b"0000_0001_0111_0000_0_0_00_0000_00000000", -- #RJMP (mode, ---, adr)  ; AR := PC
   b"0001_0100_0010_0000_0_0_00_0000_00000000", --                         ; AR := PM(adr) + AR (noflag)
   b"0000_0000_0000_0000_0_0_00_0011_00000000", --                         ; PC := AR, uPC := 0
   b"0000_0000_0000_0000_0_0_00_0101_00000000", -- #BEQ  (mode, ---, adr)  ; uPC := 0  om Z=0
   b"0000_0000_0000_0000_0_0_00_1010_00110011", --                         ; uPC := 51 om Z=1
   b"0000_0000_0000_0000_0_0_00_1010_00000000", -- #BNE  (mode, ---, adr)  ; uPC := 0  om Z=1
   b"0000_0000_0000_0000_0_0_00_0101_00110010", --                         ; uPC := 51(50) om Z=0
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_1000_0110_0_0_00_0011_00000000", -- #RIV  (----, grx, ---)  ; GrX := InputVec, uPC := 0
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --

   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000", --
   b"0000_0000_0000_0000_0_0_00_0000_00000000"  --
   );

signal u_mem : u_mem_t := u_mem_c;

begin  -- Behavioral
  uData <= u_mem(to_integer(uAddr));

end Behavioral;
